module FBCV_FORCE
(
input [15:0] IR_Prime_16,
output [15:0] FBC_V
);

assign FBC_V[11:0] = IR_Prime_16[11:0];
assign FBC_V[15:12] = 0;

endmodule
