module bit32
(
	input [15:0] valueX, //the value of X
	output [15:0] buff //output of buffer
);
assign buff[0] = 0;
assign buff[1] = 0;
assign buff[2] = valueX[0];
assign buff[3] = valueX[1];
assign buff[4] = valueX[2];
assign buff[5] = valueX[3];
assign buff[6] = valueX[4];
assign buff[7] = valueX[5];
assign buff[8] = valueX[6];
assign buff[9] = valueX[7];
assign buff[10] = valueX[8];
assign buff[11] = valueX[9];
assign buff[12] = valueX[10];
assign buff[13] = valueX[11];
assign buff[14] = valueX[12];
assign buff[15] = valueX[13];

endmodule
